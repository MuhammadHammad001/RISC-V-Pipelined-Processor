module mux4x1(inp1, inp2, inp3, sel, out);
    input   logic [31:0]    inp1;
    input   logic [31:0]    inp2;
    input   logic [31:0]    inp3;
    input   logic [1:0]     sel ;
    output  logic [31:0]    out ;


endmodule