module fetch();

endmodule