module PipelinedProcessor(clk, rst_n);
    //TODO: Complete this after adding Floating Point Unit Support.

endmodule
